// osscilator.v

// Generated using ACDS version 23.1 991

`timescale 1 ps / 1 ps
module osscilator (
		output wire  clkout, // clkout.clk
		input  wire  oscena  // oscena.oscena
	);

	altera_int_osc int_osc_0 (
		.oscena (oscena), // oscena.oscena
		.clkout (clkout)  // clkout.clk
	);

endmodule
