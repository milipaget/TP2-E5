
module osscilator (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
